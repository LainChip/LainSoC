module axi2hpi (
    input soc_clk,
    input reset,


    AXI_BUS.Slave   slv
);

endmodule